.SUBCKT irlru8726 1 2 3
* SPICE3 MODEL WITH THERMAL RC NETWORK
* Model generated on May 15, 09
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=2.60152 LAMBDA=0.00253956 KP=162.96
+CGSO=1.9685e-05 CGDO=7.85118e-07
RS 8 3 0.0022798
D1 3 1 MD
.MODEL MD D IS=1.92955e-08 RS=0.00264461 N=1.25557 BV=30
+IBV=0.00025 EG=1 XTI=2.90479 TT=1e-07
+CJO=7.19887e-10 VJ=5 M=0.731211 FC=0.5
RDS 3 1 4e+07
RD 9 1 0.0001
RG 2 7 5.695
D2 4 5 MD1
.MODEL MD1 D IS=1e-32 N=50
+CJO=3.58396e-10 VJ=0.5 M=0.3 FC=1e-08
D3 0 5 MD2
.MODEL MD2 D IS=1e-10 N=0.4 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 1.19743e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
.MODEL MD3 D IS=1e-10 N=0.4
.ENDS irlru8726

