.SUBCKT irlp3034pbf 1 2 3
* 
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=2.39395 LAMBDA=0.0267635 KP=1000
+CGSO=9.74129e-05 CGDO=3.44361e-06
RS 8 3 0.000768834
D1 3 1 MD
.MODEL MD D IS=2.95015e-08 RS=0.00113605 N=1.14564 BV=40
+IBV=0.00025 EG=1 XTI=2.76895 TT=1e-07
+CJO=8.32027e-09 VJ=0.5 M=0.521029 FC=0.5
RDS 3 1 1e+07
RD 9 1 0.000560504
RG 2 7 6.8142
D2 4 5 MD1
.MODEL MD1 D IS=1e-32 N=50
+CJO=3.00067e-09 VJ=0.500357 M=0.412917 FC=1e-08
D3 0 5 MD2
.MODEL MD2 D IS=1e-10 N=0.40041 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 9.8109e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
.MODEL MD3 D IS=1e-10 N=0.40041
.ENDS irlp3034pbf


