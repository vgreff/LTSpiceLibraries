.SUBCKT irlb4030pbf 1 2 3
* Model generated on Oct 11, 18
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=2.38692 LAMBDA=0.0320894 KP=534.97
+CGSO=0.00011116 CGDO=2.00849e-06
RS 8 3 0.000768666
D1 3 1 MD
.MODEL MD D IS=3.30329e-09 RS=0.00156078 N=1.06517 BV=100
+IBV=0.00025 EG=1.00577 XTI=2.98727 TT=1e-07
+CJO=7.90871e-09 VJ=0.5 M=0.651347 FC=0.5
RDS 3 1 5e+07
RD 9 1 0.00220278
RG 2 7 9.76611
D2 4 5 MD1
.MODEL MD1 D IS=1e-32 N=50
+CJO=3.82909e-09 VJ=0.500314 M=0.837977 FC=1e-08
D3 0 5 MD2
.MODEL MD2 D IS=1e-10 N=0.414203 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 3.82909e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
.MODEL MD3 D IS=1e-10 N=0.414203
.ENDS irlb4030pbf
