* K544UD2A OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* 
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | | FCORRECTION PIN 1
*                | | | | | | FCORRECTION PIN 8
*                | | | | | | |
.SUBCKT 544UD2A   In+ In- V+ V- OUT FC1 FC8
Q2 N005 N001 V+ PN
Q3 N001 N001 V+ PN
Q12 N001 N001 V+ PN
Q17 N006 N001 V+ PN
Q4 N012 N005 N001 PN
Q13 N013 N006 N001 PN
Q5 N016 N015 N012 PN
Q14 N017 N015 N013 PN
Q8 N010 N010 N015 0 NP
J1 N005 In- N021 NJ
J18 N006 In+ N021 NJ
Q15 N017 N027 N035 NP
Q16 N035 N034 N042 NP
Q9 N024 N016 N027 NP
Q6 N016 N027 N034 NP
Q7 N034 N034 N041 NP
Q10 N031 N031 N040 NP
Q11 N040 N040 V- NP
Q20 N037 N036 N044 NP
Q19 N021 N029 N037 NP
Q21 N021 N026 N029 NP
Q24 N026 N029 N036 NP
Q25 N036 N036 N045 NP
Q23 N023 N014 N026 NP
R1 N044 V- 230
R2 N045 V- 430
R3 N014 N023 110
R4 N010 N006 750
R5 N005 N010 750
R6 N009 N005 4k
R7 N027 N031 30k
R8 N042 V- 240
R9 N041 V- 240
Q26 N008 N002 V+ PN
Q22 N014 N008 N002 PN
Q27 N008 N008 N015 NP
R10 V+ N002 1k6
R11 N006 N007 1k
R12 FC1 N006 200
Q28 N019 N023 N026 NP
R13 N015 N019 27k
R14 V+ N003 40k
D1 FC8 N003 DX
R15 FC8 N011 40k
D2 N015 N011 DX
C1 FC8 N017 15p 
J34 V+ N017 N018 NJ
Q38 V+ N018 N020 NP 
Q33 N007 N004 V+ PN
R16 V+ N004 36
R19 N043 V- 36
Q41 N004 N020 N022 NP 1
R20 N022 OUT 36
R21 OUT N028 36
Q42 N043 N030 N028 PN 3
Q39 N020 N020 N025 NP
Q35 N020 N025 N030 NP
R17 N025 N030 40k
Q40 N036 N043 V- NP
Q37 N039 N036 N047 NP
R18 N047 V-  240
Q31 N038 N036 N046 NP
R22 N046 V- 560
Q29 N032 N032 N036 NP
R23 N029 N032 6k6
Q30 N018 N029 N038 NP
Q36 N030 N033 N039 NP
Q32 V- N036 N033 PN 
R24 N019 N033 18k
D3 N017 N024 DX
CKP3 IN+ 0 {CKP} 
CKP2 IN-  0 {CKP} 
CKP1 FC1 0 {CKP}
CKP8 FC8 0 {CKP} 
CKP5 N009 0 {CKP} 
.param CKP=1p
.model NJ NJF(VTO=-0.9 BETA=1.6m LAMBDA=0.02 RD=36 RS=30 IS=1f CGD=1p CGS=1p PB=0.5 B=1.2 KF=1E-16 AF=1.4 FC=0.5 isr=20p)
.model NP NPN(BF=120 Cje=.25p Cjc=0.25p  mjc=0.5 VAF=80 tf=50p  VTF=5  rb=150   Re=10 Rc=20 ikf=10m Xcjc=0.1 cjs=5p mjs=0.5 is=0.1f  VJE=0.9 )
.model PN PNP (BF=25 Cje=.25p Cjc=0.25p mjc=0.5  VAF=40 tf=100p  VTF=5 rb=150  cjs=1p mjs=0.5 Re=10  rc=10 Ikf=3.3m is=0.1f VJE=0.9)
.model DX D(Is=2.52n  Rs=1 N=1.752 Cjo=0.4p M=.4 Tt=20n)
.ends K544UD2A

