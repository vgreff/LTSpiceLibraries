.SUBCKT auirgdc0250 1 2 3
*Model generated on Nov 29, 12
* MODEL FORMAT: SPICE3
*Symmetry IGBT Model (Version 1.0)
*External Node Designations
*Node 1 -> a
*Node 2 -> g
*Node 3 -> k
M1 9 6 8 8 MSUB L=100u W=100u
.MODEL MSUB NMOS LEVEL=1
+VTO=6.1702 KP=0.912047 LAMBDA=0 CGSO=3.85236e-05
RD 7 9 0.000999241
RS 4 8 0.00127093
Q1 4 7 1 QSUB OFF
.MODEL QSUB PNP
+IS=1e-17 BF=23.301 NF=0.85 VAF=448.285
+IKF=2835.09 ISE=1.04627e-11 NE=1.63177 BR=4.2428
+NR=0.75 VAR=108.347 IKR=1020.91 ISC=9.99594e-12
+NC=1.99441 RB=0.146259 IRB=101.227 RBM=0.00946154
+RE=0.0012401 RC=0.000979748 XTB=0 XTI=3.14402
+EG=1.2 CJC=1.55681e-09 VJC=0.4 MJC=0.557644
+CJE=3.11362e-08 VJE=0.4 MJE=0.9 TF=5.71019e-08
RDS 7 4 1e8
RER 4 3 0.0005
RG 6 2 5.31551
RL 10 11 1
D2 12 11 DCAP
.MODEL DCAP D IS=1e-32 N=50
+CJO=1.65502e-10 VJ=1.25111 M=0.495918 FC=0.157043
D3 0 11 DL
.MODEL DL D IS=1e-10 N=0.4
VFI2 12 0 0
FI2 6 7 VFI2 -1
EV 10 0 7 6 1
CAP 10 13 6.24213e-09
RCAP 10 14 1
D4 0 14 DL
VFI1 13 14 0
FI1 6 7 VFI1 -1
.ENDS auirgdc0250


