.SUBCKT IRF9610 1 2 3
* Model generated on Sep 8, 97
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
* RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM PMOS LEVEL=1 IS=1e-32
+VTO=-3.56894 LAMBDA=2.66635e-07 KP=0.534832
+CGSO=1.5436e-06 CGDO=1.53305e-08
RS 8 3 0.221689
D1 1 3 MD
.MODEL MD D IS=5e-09 RS=0.01 N=1 BV=300
+IBV=10 EG=1.11 XTI=3 TT=6.6752e-10
+CJO=1.54088e-10 VJ=2.99942 M=0.80296 FC=0.5
RDS 3 1 1e+06
RD 9 1 1.8028
RG 2 7 2.18034
D2 5 4 MD1
* Default values used in MD1:
* RS=0 EG=1.11 XTI=3.0 TT=0
* BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=1.92701e-10 VJ=0.856605 M=0.783168 FC=1e-08
D3 5 0 MD2
* Default values used in MD2:
* EG=1.11 XTI=3.0 TT=0 CJO=0
* BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.4 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 2.99982e-10
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 6 0 MD3
* Default values used in MD3:
* EG=1.11 XTI=3.0 TT=0 CJO=0
* RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.4
.ENDS irf9610
