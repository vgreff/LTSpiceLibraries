

* LM358LV - Rev. A
* Created by Paul Goedeke; June 06, 2018
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2018 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt LM358LV IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************


I_OS        ESDn MID 7P
I_B         31 MID 10P
V_GRp       56 MID 195
V_GRn       57 MID -195
V_ISCp      50 MID 40
V_ISCn      51 MID -40
V_ORn       39 VCLP -1.45
V11         55 38 0
V_ORp       37 VCLP 1.5
V12         54 36 0
V4          27 OUT 0
VCM_MIN     77 VEE_B -100M
VCM_MAX     78 VCC_B -1.5
I_Q         VCC VEE 125U
V_OS        85 31 2.99M
C30         21 22 15.92U  
R85         22 MID R_NOISELESS 30K 
R84         22 21 R_NOISELESS 10K 
R83         21 MID R_NOISELESS 1 
GVCCS10     24 MID 23 MID  -1
C29         25 MID 19.89F  
R82         23 25 R_NOISELESS 10K 
R81         23 26 R_NOISELESS 70K 
R80         26 MID R_NOISELESS 1 
GVCCS9      26 MID 22 MID  -3.8
GVCCS4      21 MID CL_CLAMP 27  -87
R79         28 MID R_NOISELESS 1 
XU1         29 MID MID 28 VCCS_LIM_ZO_0
R78         29 MID R_NOISELESS 101 
C22         29 24 15.92F 
R65         29 24 R_NOISELESS 10K 
R64         24 MID R_NOISELESS 1 
R63         27 28 R_NOISELESS 400K 
XCLAWn      MID VIMON VEE_B 30 VCCS_LIM_CLAW-_0
Xe_n        ESDp 31 VNSE_0
Xi_nn       ESDn MID FEMT_0_0
Xi_np       MID 31 FEMT_0_0
S5          VEE ESDp VEE ESDp  S_VSWITCH_1
S4          VEE ESDn VEE ESDn  S_VSWITCH_2
S2          ESDn VCC ESDn VCC  S_VSWITCH_3
S3          ESDp VCC ESDp VCC  S_VSWITCH_4
C28         32 MID 1P 
R77         33 32 R_NOISELESS 100 
C27         34 MID 1P 
R76         35 34 R_NOISELESS 100 
R75         MID 36 R_NOISELESS 1 
GVCCS8      36 MID 37 MID  -1
R74         38 MID R_NOISELESS 1 
GVCCS7      38 MID 39 MID  -1
C25         40 MID 25F 
R69         MID 40 R_NOISELESS 1MEG 
GVCCS6      40 MID VSENSE MID  -1U
C20         CLAMP MID 151.6N 
R68         MID CLAMP R_NOISELESS 1MEG 
XVCCS_LIM_2 41 MID MID CLAMP VCCS_LIM_2_0
R44         MID 41 R_NOISELESS 1MEG 
XVCCS_LIM_1 42 43 MID 41 VCCS_LIM_1_0
Rdummy      MID 27 R_NOISELESS 40K 
R61         MID 44 R_NOISELESS 273.3609 
C16         44 45 1.1018N 
R58         45 44 R_NOISELESS 100MEG 
GVCCS2      45 MID VEE_B MID  -258.98M
R57         MID 45 R_NOISELESS 1 
R56         MID 46 R_NOISELESS 273.3609 
C15         46 47 1.1018N 
R55         47 46 R_NOISELESS 100MEG 
GVCCS1      47 MID VCC_B MID  -258.98M
R54         MID 47 R_NOISELESS 1 
R49         MID 48 R_NOISELESS 337.4K 
C14         48 49 591.7F 
R48         49 48 R_NOISELESS 100MEG 
G_adjust    49 MID ESDp MID  -44.81M
Rsrc        MID 49 R_NOISELESS 1 
XIQPos      VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQNeg      MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 2P 
XCL_AMP     50 51 VIMON MID 52 53 CLAMP_AMP_LO_0
SOR_SWp     CLAMP 54 CLAMP 54  S_VSWITCH_5
SOR_SWn     55 CLAMP 55 CLAMP  S_VSWITCH_6
XGR_AMP     56 57 58 MID 59 60 CLAMP_AMP_HI_0
R39         56 MID R_NOISELESS 1T 
R37         57 MID R_NOISELESS 1T 
R42         VSENSE 58 R_NOISELESS 1M 
C19         58 MID 1F 
R38         59 MID R_NOISELESS 1 
R36         MID 60 R_NOISELESS 1 
R40         59 61 R_NOISELESS 1M 
R41         60 62 R_NOISELESS 1M 
C17         61 MID 1F 
C18         MID 62 1F 
XGR_SRC     61 62 CLAMP MID VCCS_LIM_GR_0
R21         52 MID R_NOISELESS 1 
R20         MID 53 R_NOISELESS 1 
R29         52 63 R_NOISELESS 1M 
R30         53 64 R_NOISELESS 1M 
C9          63 MID 1F 
C8          MID 64 1F 
XCL_SRC     63 64 CL_CLAMP MID VCCS_LIM_4_0
R22         50 MID R_NOISELESS 1T 
R19         MID 51 R_NOISELESS 1T 
XCLAWp      VIMON MID 65 VCC_B VCCS_LIM_CLAW+_0
R12         65 VCC_B R_NOISELESS 1K 
R16         65 66 R_NOISELESS 1M 
R13         VEE_B 30 R_NOISELESS 1K 
R17         67 30 R_NOISELESS 1M 
C6          67 MID 1F 
C5          MID 66 1F 
G2          VCC_CLP MID 66 MID  -1M
R15         VCC_CLP MID R_NOISELESS 1K 
G3          VEE_CLP MID 67 MID  -1M
R14         MID VEE_CLP R_NOISELESS 1K 
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 68 69 CLAMP_AMP_LO_0
R26         VCC_CLP MID R_NOISELESS 1T 
R23         VEE_CLP MID R_NOISELESS 1T 
R25         68 MID R_NOISELESS 1 
R24         MID 69 R_NOISELESS 1 
R27         68 70 R_NOISELESS 1M 
R28         69 71 R_NOISELESS 1M 
C11         70 MID 1F 
C10         MID 71 1F 
XCLAW_SRC   70 71 CLAW_CLAMP MID VCCS_LIM_3_0
H2          35 MID V11 -1
H3          33 MID V12 1
C12         SW_OL MID 100P 
R32         72 SW_OL R_NOISELESS 100 
R31         72 MID R_NOISELESS 1 
XOL_SENSE   MID 72 34 32 OL_SENSE_0
S1          21 22 SW_OL MID  S_VSWITCH_7
H1          73 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_8
S6          OUT VCC OUT VCC  S_VSWITCH_9
R11         MID 74 R_NOISELESS 1T 
R18         74 VOUT_S R_NOISELESS 100 
C7          VOUT_S MID 1P 
E5          74 MID OUT MID  1
C13         VIMON MID 1N 
R33         73 VIMON R_NOISELESS 100 
R10         MID 73 R_NOISELESS 1T 
R47         75 VCLP R_NOISELESS 100 
C24         VCLP MID 100P 
E4          75 MID CL_CLAMP MID  1
R46         MID CL_CLAMP R_NOISELESS 1K 
G9          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP R_NOISELESS 1K 
G8          CLAW_CLAMP MID 40 MID  -1M
R43         MID VSENSE R_NOISELESS 1K 
G15         VSENSE MID CLAMP MID  -1M
C4          42 MID 1F 
R9          42 76 R_NOISELESS 1M 
R7          MID 77 R_NOISELESS 1T 
R6          78 MID R_NOISELESS 1T 
R8          MID 76 R_NOISELESS 1 
XVCM_CLAMP  79 MID 76 MID 78 77 VCCS_EXT_LIM_0
E1          MID 0 80 0  1
R89         VEE_B 0 R_NOISELESS 1 
R5          81 VEE_B R_NOISELESS 1M 
C3          81 0 1F 
R60         80 81 R_NOISELESS 1MEG 
C1          80 0 1 
R3          80 0 R_NOISELESS 1T 
R59         82 80 R_NOISELESS 1MEG 
C2          82 0 1F 
R4          VCC_B 82 R_NOISELESS 1M 
R88         VCC_B 0 R_NOISELESS 1 
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R_PSR       83 79 R_NOISELESS 1K 
G_PSR       79 83 46 44  -1M
R2          43 ESDn R_NOISELESS 1M 
R1          83 84 R_NOISELESS 1M 
R_CMR       85 84 R_NOISELESS 1K 
G_CMR       84 85 48 MID  -1M
C_CMn       ESDn MID 5.5P 
C_CMp       MID ESDp 5.5P 
R53         ESDn MID R_NOISELESS 1T 
R52         MID ESDp R_NOISELESS 1T 
R35         IN- ESDn R_NOISELESS 10M 
R34         IN+ ESDp R_NOISELESS 10M 

.MODEL S_VSWITCH_1 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_2 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_3 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_5 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_6 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_7 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_8 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_9 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)

*$
*
.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 100
.PARAM IPOS = 32E3
.PARAM INEG = -32E3
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAW-_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(00.0000, 0.00001)
+(14.0000, 0.000379)
+(28.0000, 0.000877)
+(37.3333, 0.001382)
+(37.8000, 0.00142)
+(38.7333, 0.001493)
+(39.6667, 0.001583)
+(40.6000, 0.001703)
+(41.5333, 0.00191)
+(42.0000, 0.00204)
.ENDS VCCS_LIM_CLAW-_0 
*


.SUBCKT VNSE_0  1 2
.PARAM FLW=10
.PARAM NLF=115
.PARAM NVR=27
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
*


.SUBCKT FEMT_0_0   1 2
.PARAM FLWF=0.001
.PARAM NLFF=23
.PARAM NVRF=23
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*


.SUBCKT VCCS_LIM_2_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 11.15E-3
.PARAM IPOS = 0.263
.PARAM INEG = -0.263
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.55
.PARAM INEG = -0.55
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 1.122
.PARAM INEG = -1.122
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAW+_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(00.00, 0.000010)
+(13.67, 0.0003467)
+(27.33, 0.0007994)
+(36.44, 0.001309)
+(36.90, 0.001351)
+(37.81, 0.001455)
+(38.72, 0.001600)
+(39.63, 0.001812)
+(40.54, 0.002117)
+(41.00, 0.002292)
.ENDS VCCS_LIM_CLAW+_0 
*


.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.47
.PARAM INEG = -0.47
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
.ENDS LM358LV
*

* LMX58B_LM2904B - Rev. A
* Created by Paul Goedeke; November 19, 2018
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2018 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.SUBCKT LMX58B_LM2904B  IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************


I_OS        ESDn MID -9.5N
I_B         37 MID -10N
V_GRp       57 MID 180
V_GRn       58 MID -180
V_ISCp      51 MID 40
V_ISCn      52 MID -40
V_ORn       45 VCLP -1.2
V11         56 44 0
V_ORp       43 VCLP 1.2
V12         55 42 0
V4          33 OUT 0
VCM_MIN     79 VEE_B 0
VCM_MAX     80 VCC_B -1.5
I_Q         VCC VEE 300U
V_OS        86 37 264U
R57         MID 22 R_NOISELESS 1K 
C16         22 23 1.592P 
R51         23 22 R_NOISELESS 100MEG 
GVCCS2      23 MID VEE_B MID  -100M
R50         MID 23 R_NOISELESS 1 
XU3         VCC_B VEE_B 24 25 26 27 MID PHASEREV_0
XU1         VIMON MID CRS CRS_DIST_0
C21         28 29 313.8N  
C22         30 31 636.6F  
R70         31 MID R_NOISELESS 2.5 
R67         31 30 R_NOISELESS 10K 
R66         30 MID R_NOISELESS 1 
XU2         31 MID MID 32 VCCS_LIM_ZO_0
GVCCS4      30 MID 29 MID  -4.3
R65         29 MID R_NOISELESS 3.03K 
R64         29 28 R_NOISELESS 10K 
R63         28 MID R_NOISELESS 1 
GVCCS3      28 MID CL_CLAMP 33  -90
R62         32 MID R_NOISELESS 1 
C29         34 MID 47F 
R78         MID 34 R_NOISELESS 1MEG 
GVCCS9      34 MID 35 MID  -1U
XU5         36 MID MID CLAMP CRS MID VCCS_LIM_2_EN_0
C28         38 MID 1P 
R77         39 38 R_NOISELESS 100 
C27         40 MID 1P 
R76         41 40 R_NOISELESS 100 
R75         MID 42 R_NOISELESS 1 
GVCCS8      42 MID 43 MID  -1
R74         44 MID R_NOISELESS 1 
GVCCS7      44 MID 45 MID  -1
Xi_nn       ESDn MID FEMT_0
Xi_np       MID 37 FEMT_0
Xe_n        ESDp 37 VNSE_0
C25         35 MID 47F 
R69         MID 35 R_NOISELESS 1MEG 
GVCCS6      35 MID VSENSE MID  -1U
C20         CLAMP MID 9N 
R68         MID CLAMP R_NOISELESS 1MEG 
R44         MID 36 R_NOISELESS 1MEG 
XVCCS_LIM_1 46 27 MID 36 VCCS_LIM_1_0
Rdummy      MID 33 R_NOISELESS 25K 
Rx          33 32 R_NOISELESS 250K 
R56         MID 47 R_NOISELESS 1K 
C15         47 48 1.592P 
R55         48 47 R_NOISELESS 100MEG 
GVCCS1      48 MID VCC_B MID  -100M
R54         MID 48 R_NOISELESS 1 
R49         MID 49 R_NOISELESS 4.616K 
C14         49 50 26.53P 
R48         50 49 R_NOISELESS 100MEG 
G_adjust    50 MID ESDp MID  -685.2M
Rsrc        MID 50 R_NOISELESS 1 
XIQPos      VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQNeg      MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 1P 
XCL_AMP     51 52 VIMON MID 53 54 CLAMP_AMP_LO_0
SOR_SWp     CLAMP 55 CLAMP 55  S_VSWITCH_1
SOR_SWn     56 CLAMP 56 CLAMP  S_VSWITCH_2
XGR_AMP     57 58 59 MID 60 61 CLAMP_AMP_HI_0
R39         57 MID R_NOISELESS 1T 
R37         58 MID R_NOISELESS 1T 
R42         VSENSE 59 R_NOISELESS 1M 
C19         59 MID 1F 
R38         60 MID R_NOISELESS 1 
R36         MID 61 R_NOISELESS 1 
R40         60 62 R_NOISELESS 1M 
R41         61 63 R_NOISELESS 1M 
C17         62 MID 1F 
C18         MID 63 1F 
XGR_SRC     62 63 CLAMP MID VCCS_LIM_GR_0
R21         53 MID R_NOISELESS 1 
R20         MID 54 R_NOISELESS 1 
R29         53 64 R_NOISELESS 1M 
R30         54 65 R_NOISELESS 1M 
C9          64 MID 1F 
C8          MID 65 1F 
XCL_SRC     64 65 CL_CLAMP MID VCCS_LIM_4_0
R22         51 MID R_NOISELESS 1T 
R19         MID 52 R_NOISELESS 1T 
XCLAWp      VIMON MID 66 VCC_B VCCS_LIM_CLAW+_0
XCLAWn      MID VIMON VEE_B 67 VCCS_LIM_CLAW-_0
R12         66 VCC_B R_NOISELESS 1K 
R16         66 68 R_NOISELESS 1M 
R13         VEE_B 67 R_NOISELESS 1K 
R17         69 67 R_NOISELESS 1M 
C6          69 MID 1F 
C5          MID 68 1F 
G2          VCC_CLP MID 68 MID  -1M
R15         VCC_CLP MID R_NOISELESS 1K 
G3          VEE_CLP MID 69 MID  -1M
R14         MID VEE_CLP R_NOISELESS 1K 
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 70 71 CLAMP_AMP_LO_0
R26         VCC_CLP MID R_NOISELESS 1T 
R23         VEE_CLP MID R_NOISELESS 1T 
R25         70 MID R_NOISELESS 1 
R24         MID 71 R_NOISELESS 1 
R27         70 72 R_NOISELESS 1M 
R28         71 73 R_NOISELESS 1M 
C11         72 MID 1F 
C10         MID 73 1F 
XCLAW_SRC   72 73 CLAW_CLAMP MID VCCS_LIM_3_0
H2          41 MID V11 -1
H3          39 MID V12 1
C12         SW_OL MID 100P 
R32         74 SW_OL R_NOISELESS 100 
R31         74 MID R_NOISELESS 1 
XOL_SENSE   MID 74 40 38 OL_SENSE_0
S1          28 29 SW_OL MID  S_VSWITCH_3
H1          75 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_4
S6          OUT VCC OUT VCC  S_VSWITCH_5
R11         MID 76 R_NOISELESS 1T 
R18         76 VOUT_S R_NOISELESS 100 
C7          VOUT_S MID 10P 
E5          76 MID OUT MID  1
C13         VIMON MID 10P 
R33         75 VIMON R_NOISELESS 100 
R10         MID 75 R_NOISELESS 1T 
R47         77 VCLP R_NOISELESS 100 
C24         VCLP MID 100P 
E4          77 MID CL_CLAMP MID  1
R46         MID CL_CLAMP R_NOISELESS 1K 
G9          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP R_NOISELESS 1K 
G8          CLAW_CLAMP MID 34 MID  -1M
R43         MID VSENSE R_NOISELESS 1K 
G15         VSENSE MID CLAMP MID  -1M
C4          46 MID 1F 
R9          46 78 R_NOISELESS 1M 
R7          MID 79 R_NOISELESS 1T 
R6          80 MID R_NOISELESS 1T 
R8          MID 78 R_NOISELESS 1 
XVCM_CLAMP  26 MID 78 MID 80 79 VCCS_EXT_LIM_0
E1          MID 0 81 0  1
R89         VEE_B 0 R_NOISELESS 1 
R5          82 VEE_B R_NOISELESS 1M 
C3          82 0 1F 
R60         81 82 R_NOISELESS 1MEG 
C1          81 0 1 
R3          81 0 R_NOISELESS 1T 
R59         83 81 R_NOISELESS 1MEG 
C2          83 0 1F 
R4          VCC_B 83 R_NOISELESS 1M 
R88         VCC_B 0 R_NOISELESS 1 
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R_PSR       84 24 R_NOISELESS 1K 
G_PSR       24 84 47 22  -1M
R2          25 ESDn R_NOISELESS 1M 
R1          84 85 R_NOISELESS 1M 
R_CMR       86 85 R_NOISELESS 1K 
G_CMR       85 86 49 MID  -1M
C_CMn       ESDn MID 2P 
C_CMp       MID ESDp 2P 
R53         ESDn MID R_NOISELESS 1T 
R52         MID ESDp R_NOISELESS 1T 
R35         IN- ESDn R_NOISELESS 10M 
R34         IN+ ESDp R_NOISELESS 10M 

.MODEL S_VSWITCH_1 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_2 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_3 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_5 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
*
*$
*
.SUBCKT PHASEREV_0  VCC VEE VIN+ VIN- VOUT+ VOUT- MID
E1 VOUT+ MID VALUE={IF(V(VIN+,MID)<V(VEE,MID)-0.3,V(VCC,MID),V(VIN+,MID))}
E2 VOUT- MID VALUE={IF(V(VIN-,MID)<V(VEE,MID)-0.3,V(VCC,MID),V(VIN-,MID))}
.ENDS
*


.SUBCKT CRS_DIST_0  VIMON MID OUT
V1 VREF MID -40M
ESHF VSHF MID VIMON VREF 1
GZC MID ZC VALUE = {SGN(V(VSHF,MID))}
R1 ZC MID 1
C1 ZC MID 2U
GCR MID OUT VALUE = {IF((ABS(V(ZC,MID))<=0.9),0,1)}
R2 OUT MID 1
.ENDS
*


.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 4E3
.PARAM IPOS = 1E6
.PARAM INEG = -1E6
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_2_EN_0  VC+ VC- IOUT+ IOUT- EN MID
.PARAM GAIN = 8.4E-4
.PARAM IPOS = 0.0048
.PARAM INEG = -0.0048
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(EN,MID)*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT FEMT_0  1 2
.PARAM FLWF=1E-3
.PARAM NLFF=500
.PARAM NVRF=500
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*


.SUBCKT VNSE_0  1 2
.PARAM FLW=10
.PARAM NLF=80
.PARAM NVR=35
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
*


.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.013
.PARAM INEG = -0.013
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 1.04
.PARAM INEG = -1.04
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAW+_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 1.17E-03)
+(0.0046251, 1.17E-3)
+(0.15716, 1.21E-3)
+(1.3309, 1.28E-3)
+(35.075, 2.12E-3)
+(35.680, 2.55E-3)
+(36.033, 2.84E-3)
+(37.416, 7.97E-3)
.ENDS
*


.SUBCKT VCCS_LIM_CLAW-_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0.010, 2.50E-5)
+(0.070, 2.50E-5)
+(0.090, 5.80E-4)
+(0.100, 6.06E-4)
+(0.760, 7.14E-4) 
+(1.440, 7.62E-4)
+(8.000, 1.10E-3)
+(13.60, 1.55E-3)
+(15.45, 1.75E-3)
+(17.26, 2.15E-3)
+(18.87, 2.94E-3)
+(21.58, 4.50E-3)
+(25.53, 1.02E-2)
.ENDS
*



.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.435
.PARAM INEG = -0.435
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
.ENDS LMX58B_LM2904B
*

* LM358BTI - Rev. A
* Created by Paul Goedeke; November 19, 2018
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2018 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt LM358BTI  IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************


I_OS        ESDn MID -9.5N
I_B         37 MID -10N
V_GRp       57 MID 180
V_GRn       58 MID -180
V_ISCp      51 MID 40
V_ISCn      52 MID -40
V_ORn       45 VCLP -1.2
V11         56 44 0
V_ORp       43 VCLP 1.2
V12         55 42 0
V4          33 OUT 0
VCM_MIN     79 VEE_B 0
VCM_MAX     80 VCC_B -1.5
I_Q         VCC VEE 300U
V_OS        86 37 264U
R57         MID 22 R_NOISELESS 1K 
C16         22 23 1.592P 
R51         23 22 R_NOISELESS 100MEG 
GVCCS2      23 MID VEE_B MID  -100M
R50         MID 23 R_NOISELESS 1 
XU3         VCC_B VEE_B 24 25 26 27 MID PHASEREV_0
XU1         VIMON MID CRS CRS_DIST_0
C21         28 29 313.8N  
C22         30 31 636.6F  
R70         31 MID R_NOISELESS 2.5 
R67         31 30 R_NOISELESS 10K 
R66         30 MID R_NOISELESS 1 
XU2         31 MID MID 32 VCCS_LIM_ZO_0
GVCCS4      30 MID 29 MID  -4.3
R65         29 MID R_NOISELESS 3.03K 
R64         29 28 R_NOISELESS 10K 
R63         28 MID R_NOISELESS 1 
GVCCS3      28 MID CL_CLAMP 33  -90
R62         32 MID R_NOISELESS 1 
C29         34 MID 47F 
R78         MID 34 R_NOISELESS 1MEG 
GVCCS9      34 MID 35 MID  -1U
XU5         36 MID MID CLAMP CRS MID VCCS_LIM_2_EN_0
C28         38 MID 1P 
R77         39 38 R_NOISELESS 100 
C27         40 MID 1P 
R76         41 40 R_NOISELESS 100 
R75         MID 42 R_NOISELESS 1 
GVCCS8      42 MID 43 MID  -1
R74         44 MID R_NOISELESS 1 
GVCCS7      44 MID 45 MID  -1
Xi_nn       ESDn MID FEMT_0
Xi_np       MID 37 FEMT_0
Xe_n        ESDp 37 VNSE_0
C25         35 MID 47F 
R69         MID 35 R_NOISELESS 1MEG 
GVCCS6      35 MID VSENSE MID  -1U
C20         CLAMP MID 9N 
R68         MID CLAMP R_NOISELESS 1MEG 
R44         MID 36 R_NOISELESS 1MEG 
XVCCS_LIM_1 46 27 MID 36 VCCS_LIM_1_0
Rdummy      MID 33 R_NOISELESS 25K 
Rx          33 32 R_NOISELESS 250K 
R56         MID 47 R_NOISELESS 1K 
C15         47 48 1.592P 
R55         48 47 R_NOISELESS 100MEG 
GVCCS1      48 MID VCC_B MID  -100M
R54         MID 48 R_NOISELESS 1 
R49         MID 49 R_NOISELESS 4.616K 
C14         49 50 26.53P 
R48         50 49 R_NOISELESS 100MEG 
G_adjust    50 MID ESDp MID  -685.2M
Rsrc        MID 50 R_NOISELESS 1 
XIQPos      VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQNeg      MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 1P 
XCL_AMP     51 52 VIMON MID 53 54 CLAMP_AMP_LO_0
SOR_SWp     CLAMP 55 CLAMP 55  S_VSWITCH_1
SOR_SWn     56 CLAMP 56 CLAMP  S_VSWITCH_2
XGR_AMP     57 58 59 MID 60 61 CLAMP_AMP_HI_0
R39         57 MID R_NOISELESS 1T 
R37         58 MID R_NOISELESS 1T 
R42         VSENSE 59 R_NOISELESS 1M 
C19         59 MID 1F 
R38         60 MID R_NOISELESS 1 
R36         MID 61 R_NOISELESS 1 
R40         60 62 R_NOISELESS 1M 
R41         61 63 R_NOISELESS 1M 
C17         62 MID 1F 
C18         MID 63 1F 
XGR_SRC     62 63 CLAMP MID VCCS_LIM_GR_0
R21         53 MID R_NOISELESS 1 
R20         MID 54 R_NOISELESS 1 
R29         53 64 R_NOISELESS 1M 
R30         54 65 R_NOISELESS 1M 
C9          64 MID 1F 
C8          MID 65 1F 
XCL_SRC     64 65 CL_CLAMP MID VCCS_LIM_4_0
R22         51 MID R_NOISELESS 1T 
R19         MID 52 R_NOISELESS 1T 
XCLAWp      VIMON MID 66 VCC_B VCCS_LIM_CLAW+_0
XCLAWn      MID VIMON VEE_B 67 VCCS_LIM_CLAW-_0
R12         66 VCC_B R_NOISELESS 1K 
R16         66 68 R_NOISELESS 1M 
R13         VEE_B 67 R_NOISELESS 1K 
R17         69 67 R_NOISELESS 1M 
C6          69 MID 1F 
C5          MID 68 1F 
G2          VCC_CLP MID 68 MID  -1M
R15         VCC_CLP MID R_NOISELESS 1K 
G3          VEE_CLP MID 69 MID  -1M
R14         MID VEE_CLP R_NOISELESS 1K 
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 70 71 CLAMP_AMP_LO_0
R26         VCC_CLP MID R_NOISELESS 1T 
R23         VEE_CLP MID R_NOISELESS 1T 
R25         70 MID R_NOISELESS 1 
R24         MID 71 R_NOISELESS 1 
R27         70 72 R_NOISELESS 1M 
R28         71 73 R_NOISELESS 1M 
C11         72 MID 1F 
C10         MID 73 1F 
XCLAW_SRC   72 73 CLAW_CLAMP MID VCCS_LIM_3_0
H2          41 MID V11 -1
H3          39 MID V12 1
C12         SW_OL MID 100P 
R32         74 SW_OL R_NOISELESS 100 
R31         74 MID R_NOISELESS 1 
XOL_SENSE   MID 74 40 38 OL_SENSE_0
S1          28 29 SW_OL MID  S_VSWITCH_3
H1          75 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_4
S6          OUT VCC OUT VCC  S_VSWITCH_5
R11         MID 76 R_NOISELESS 1T 
R18         76 VOUT_S R_NOISELESS 100 
C7          VOUT_S MID 10P 
E5          76 MID OUT MID  1
C13         VIMON MID 10P 
R33         75 VIMON R_NOISELESS 100 
R10         MID 75 R_NOISELESS 1T 
R47         77 VCLP R_NOISELESS 100 
C24         VCLP MID 100P 
E4          77 MID CL_CLAMP MID  1
R46         MID CL_CLAMP R_NOISELESS 1K 
G9          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP R_NOISELESS 1K 
G8          CLAW_CLAMP MID 34 MID  -1M
R43         MID VSENSE R_NOISELESS 1K 
G15         VSENSE MID CLAMP MID  -1M
C4          46 MID 1F 
R9          46 78 R_NOISELESS 1M 
R7          MID 79 R_NOISELESS 1T 
R6          80 MID R_NOISELESS 1T 
R8          MID 78 R_NOISELESS 1 
XVCM_CLAMP  26 MID 78 MID 80 79 VCCS_EXT_LIM_0
E1          MID 0 81 0  1
R89         VEE_B 0 R_NOISELESS 1 
R5          82 VEE_B R_NOISELESS 1M 
C3          82 0 1F 
R60         81 82 R_NOISELESS 1MEG 
C1          81 0 1 
R3          81 0 R_NOISELESS 1T 
R59         83 81 R_NOISELESS 1MEG 
C2          83 0 1F 
R4          VCC_B 83 R_NOISELESS 1M 
R88         VCC_B 0 R_NOISELESS 1 
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R_PSR       84 24 R_NOISELESS 1K 
G_PSR       24 84 47 22  -1M
R2          25 ESDn R_NOISELESS 1M 
R1          84 85 R_NOISELESS 1M 
R_CMR       86 85 R_NOISELESS 1K 
G_CMR       85 86 49 MID  -1M
C_CMn       ESDn MID 2P 
C_CMp       MID ESDp 2P 
R53         ESDn MID R_NOISELESS 1T 
R52         MID ESDp R_NOISELESS 1T 
R35         IN- ESDn R_NOISELESS 10M 
R34         IN+ ESDp R_NOISELESS 10M 

.MODEL S_VSWITCH_1 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_2 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_3 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_5 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)

*$
*
.SUBCKT PHASEREV_0  VCC VEE VIN+ VIN- VOUT+ VOUT- MID
E1 VOUT+ MID VALUE={IF(V(VIN+,MID)<V(VEE,MID)-0.3,V(VCC,MID),V(VIN+,MID))}
E2 VOUT- MID VALUE={IF(V(VIN-,MID)<V(VEE,MID)-0.3,V(VCC,MID),V(VIN-,MID))}
.ENDS
*


.SUBCKT CRS_DIST_0  VIMON MID OUT
V1 VREF MID -40M
ESHF VSHF MID VIMON VREF 1
GZC MID ZC VALUE = {SGN(V(VSHF,MID))}
R1 ZC MID 1
C1 ZC MID 2U
GCR MID OUT VALUE = {IF((ABS(V(ZC,MID))<=0.9),0,1)}
R2 OUT MID 1
.ENDS
*


.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 4E3
.PARAM IPOS = 1E6
.PARAM INEG = -1E6
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_2_EN_0  VC+ VC- IOUT+ IOUT- EN MID
.PARAM GAIN = 8.4E-4
.PARAM IPOS = 0.0048
.PARAM INEG = -0.0048
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(EN,MID)*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT FEMT_0  1 2
.PARAM FLWF=1E-3
.PARAM NLFF=500
.PARAM NVRF=500
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*


.SUBCKT VNSE_0  1 2
.PARAM FLW=10
.PARAM NLF=80
.PARAM NVR=35
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
*


.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.013
.PARAM INEG = -0.013
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 1.04
.PARAM INEG = -1.04
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAW+_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 1.17E-03)
+(0.0046251, 1.17E-3)
+(0.15716, 1.21E-3)
+(1.3309, 1.28E-3)
+(35.075, 2.12E-3)
+(35.680, 2.55E-3)
+(36.033, 2.84E-3)
+(37.416, 7.97E-3)
.ENDS
*


.SUBCKT VCCS_LIM_CLAW-_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0.010, 2.50E-5)
+(0.070, 2.50E-5)
+(0.090, 5.80E-4)
+(0.100, 6.06E-4)
+(0.760, 7.14E-4) 
+(1.440, 7.62E-4)
+(8.000, 1.10E-3)
+(13.60, 1.55E-3)
+(15.45, 1.75E-3)
+(17.26, 2.15E-3)
+(18.87, 2.94E-3)
+(21.58, 4.50E-3)
+(25.53, 1.02E-2)
.ENDS
*



.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.435
.PARAM INEG = -0.435
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
.ENDS LM358BTI
*

* LM358TI - Rev. A
* Created by Paul Goedeke; November 16, 2018
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2018 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt LM358TI  IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************


I_OS        ESDn MID -18N
I_B         37 MID -20N
V_GRp       57 MID 180
V_GRn       58 MID -180
V_ISCp      51 MID 40
V_ISCn      52 MID -40
V_ORn       45 VCLP -1.2
V11         56 44 0
V_ORp       43 VCLP 1.2
V12         55 42 0
V4          33 OUT 0
VCM_MIN     79 VEE_B 0
VCM_MAX     80 VCC_B -1.5
I_Q         VCC VEE 350U
V_OS        86 37 1.8M
R61         MID 22 R_NOISELESS 8.001K 
C16         22 23 19.89P 
R58         23 22 R_NOISELESS 100MEG 
GVCCS2      23 MID VEE_B MID  -992.9M
R57         MID 23 R_NOISELESS 1 
XU3         VCC_B VEE_B 24 25 26 27 MID PHASEREV_0
XU1         VIMON MID CRS CRS_DIST_0
C21         28 29 313.8N  
C22         30 31 636.6F  
R70         31 MID R_NOISELESS 2.5 
R67         31 30 R_NOISELESS 10K 
R66         30 MID R_NOISELESS 1 
XU2         31 MID MID 32 VCCS_LIM_ZO_0
GVCCS4      30 MID 29 MID  -4.3
R65         29 MID R_NOISELESS 3.03K 
R64         29 28 R_NOISELESS 10K 
R63         28 MID R_NOISELESS 1 
GVCCS3      28 MID CL_CLAMP 33  -90
R62         32 MID R_NOISELESS 1 
C29         34 MID 72F 
R78         MID 34 R_NOISELESS 1MEG 
GVCCS9      34 MID 35 MID  -1U
XU5         36 MID MID CLAMP CRS MID VCCS_LIM_2_EN_0
C28         38 MID 1P 
R77         39 38 R_NOISELESS 100 
C27         40 MID 1P 
R76         41 40 R_NOISELESS 100 
R75         MID 42 R_NOISELESS 1 
GVCCS8      42 MID 43 MID  -1
R74         44 MID R_NOISELESS 1 
GVCCS7      44 MID 45 MID  -1
Xi_nn       ESDn MID FEMT_0
Xi_np       MID 37 FEMT_0
Xe_n        ESDp 37 VNSE_0
C25         35 MID 72F 
R69         MID 35 R_NOISELESS 1MEG 
GVCCS6      35 MID VSENSE MID  -1U
C20         CLAMP MID 13.5N 
R68         MID CLAMP R_NOISELESS 1MEG 
R44         MID 36 R_NOISELESS 1MEG 
XVCCS_LIM_1 46 27 MID 36 VCCS_LIM_1_0
Rdummy      MID 33 R_NOISELESS 25K 
Rx          33 32 R_NOISELESS 250K 
R56         MID 47 R_NOISELESS 1K 
C15         47 48 1.592P 
R55         48 47 R_NOISELESS 100MEG 
GVCCS1      48 MID VCC_B MID  -100M
R54         MID 48 R_NOISELESS 1 
R49         MID 49 R_NOISELESS 4.616K 
C14         49 50 26.53P 
R48         50 49 R_NOISELESS 100MEG 
G_adjust    50 MID ESDp MID  -685.2M
Rsrc        MID 50 R_NOISELESS 1 
XIQPos      VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQNeg      MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 1P 
XCL_AMP     51 52 VIMON MID 53 54 CLAMP_AMP_LO_0
SOR_SWp     CLAMP 55 CLAMP 55  S_VSWITCH_1
SOR_SWn     56 CLAMP 56 CLAMP  S_VSWITCH_2
XGR_AMP     57 58 59 MID 60 61 CLAMP_AMP_HI_0
R39         57 MID R_NOISELESS 1T 
R37         58 MID R_NOISELESS 1T 
R42         VSENSE 59 R_NOISELESS 1M 
C19         59 MID 1F 
R38         60 MID R_NOISELESS 1 
R36         MID 61 R_NOISELESS 1 
R40         60 62 R_NOISELESS 1M 
R41         61 63 R_NOISELESS 1M 
C17         62 MID 1F 
C18         MID 63 1F 
XGR_SRC     62 63 CLAMP MID VCCS_LIM_GR_0
R21         53 MID R_NOISELESS 1 
R20         MID 54 R_NOISELESS 1 
R29         53 64 R_NOISELESS 1M 
R30         54 65 R_NOISELESS 1M 
C9          64 MID 1F 
C8          MID 65 1F 
XCL_SRC     64 65 CL_CLAMP MID VCCS_LIM_4_0
R22         51 MID R_NOISELESS 1T 
R19         MID 52 R_NOISELESS 1T 
XCLAWp      VIMON MID 66 VCC_B VCCS_LIM_CLAW+_0
XCLAWn      MID VIMON VEE_B 67 VCCS_LIM_CLAW-_0
R12         66 VCC_B R_NOISELESS 1K 
R16         66 68 R_NOISELESS 1M 
R13         VEE_B 67 R_NOISELESS 1K 
R17         69 67 R_NOISELESS 1M 
C6          69 MID 1F 
C5          MID 68 1F 
G2          VCC_CLP MID 68 MID  -1M
R15         VCC_CLP MID R_NOISELESS 1K 
G3          VEE_CLP MID 69 MID  -1M
R14         MID VEE_CLP R_NOISELESS 1K 
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 70 71 CLAMP_AMP_LO_0
R26         VCC_CLP MID R_NOISELESS 1T 
R23         VEE_CLP MID R_NOISELESS 1T 
R25         70 MID R_NOISELESS 1 
R24         MID 71 R_NOISELESS 1 
R27         70 72 R_NOISELESS 1M 
R28         71 73 R_NOISELESS 1M 
C11         72 MID 1F 
C10         MID 73 1F 
XCLAW_SRC   72 73 CLAW_CLAMP MID VCCS_LIM_3_0
H2          41 MID V11 -1
H3          39 MID V12 1
C12         SW_OL MID 100P 
R32         74 SW_OL R_NOISELESS 100 
R31         74 MID R_NOISELESS 1 
XOL_SENSE   MID 74 40 38 OL_SENSE_0
S1          28 29 SW_OL MID  S_VSWITCH_3
H1          75 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_4
S6          OUT VCC OUT VCC  S_VSWITCH_5
R11         MID 76 R_NOISELESS 1T 
R18         76 VOUT_S R_NOISELESS 100 
C7          VOUT_S MID 10P 
E5          76 MID OUT MID  1
C13         VIMON MID 10P 
R33         75 VIMON R_NOISELESS 100 
R10         MID 75 R_NOISELESS 1T 
R47         77 VCLP R_NOISELESS 100 
C24         VCLP MID 100P 
E4          77 MID CL_CLAMP MID  1
R46         MID CL_CLAMP R_NOISELESS 1K 
G9          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP R_NOISELESS 1K 
G8          CLAW_CLAMP MID 34 MID  -1M
R43         MID VSENSE R_NOISELESS 1K 
G15         VSENSE MID CLAMP MID  -1M
C4          46 MID 1F 
R9          46 78 R_NOISELESS 1M 
R7          MID 79 R_NOISELESS 1T 
R6          80 MID R_NOISELESS 1T 
R8          MID 78 R_NOISELESS 1 
XVCM_CLAMP  26 MID 78 MID 80 79 VCCS_EXT_LIM_0
E1          MID 0 81 0  1
R89         VEE_B 0 R_NOISELESS 1 
R5          82 VEE_B R_NOISELESS 1M 
C3          82 0 1F 
R60         81 82 R_NOISELESS 1MEG 
C1          81 0 1 
R3          81 0 R_NOISELESS 1T 
R59         83 81 R_NOISELESS 1MEG 
C2          83 0 1F 
R4          VCC_B 83 R_NOISELESS 1M 
R88         VCC_B 0 R_NOISELESS 1 
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R_PSR       84 24 R_NOISELESS 1K 
G_PSR       24 84 47 22  -1M
R2          25 ESDn R_NOISELESS 1M 
R1          84 85 R_NOISELESS 1M 
R_CMR       86 85 R_NOISELESS 1K 
G_CMR       85 86 49 MID  -1M
C_CMn       ESDn MID 2P 
C_CMp       MID ESDp 2P 
R53         ESDn MID R_NOISELESS 1T 
R52         MID ESDp R_NOISELESS 1T 
R35         IN- ESDn R_NOISELESS 10M 
R34         IN+ ESDp R_NOISELESS 10M 

.MODEL S_VSWITCH_1 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_2 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_3 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_5 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)

*$
*
.SUBCKT PHASEREV_0  VCC VEE VIN+ VIN- VOUT+ VOUT- MID
E1 VOUT+ MID VALUE={IF(V(VIN+,MID)<V(VEE,MID)-0.3,V(VCC,MID),V(VIN+,MID))}
E2 VOUT- MID VALUE={IF(V(VIN-,MID)<V(VEE,MID)-0.3,V(VCC,MID),V(VIN-,MID))}
.ENDS
*


.SUBCKT CRS_DIST_0  VIMON MID OUT
V1 VREF MID -40M
ESHF VSHF MID VIMON VREF 1
GZC MID ZC VALUE = {SGN(V(VSHF,MID))}
R1 ZC MID 1
C1 ZC MID 2U
GCR MID OUT VALUE = {IF((ABS(V(ZC,MID))<=0.9),0,1)}
R2 OUT MID 1
.ENDS
*


.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 4E3
.PARAM IPOS = 1E6
.PARAM INEG = -1E6
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_2_EN_0  VC+ VC- IOUT+ IOUT- EN MID
.PARAM GAIN = 8.4E-4
.PARAM IPOS = 0.005
.PARAM INEG = -0.005
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(EN,MID)*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT FEMT_0  1 2
.PARAM FLWF=1E-3
.PARAM NLFF=500
.PARAM NVRF=500
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*


.SUBCKT VNSE_0  1 2
.PARAM FLW=10
.PARAM NLF=80
.PARAM NVR=35
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
*


.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.013
.PARAM INEG = -0.013
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 1.04
.PARAM INEG = -1.04
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAW+_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 1.17E-03)
+(0.0046251, 1.17E-3)
+(0.15716, 1.21E-3)
+(1.3309, 1.28E-3)
+(35.075, 2.12E-3)
+(35.680, 2.55E-3)
+(36.033, 2.84E-3)
+(37.416, 7.97E-3)
.ENDS
*


.SUBCKT VCCS_LIM_CLAW-_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0.010, 2.50E-5)
+(0.070, 2.50E-5)
+(0.090, 5.80E-4)
+(0.100, 6.06E-4)
+(0.760, 7.14E-4) 
+(1.440, 7.62E-4)
+(8.000, 1.10E-3)
+(13.60, 1.55E-3)
+(15.45, 1.75E-3)
+(17.26, 2.15E-3)
+(18.87, 2.94E-3)
+(21.58, 4.50E-3)
+(25.53, 1.02E-2)
.ENDS
*



.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.435
.PARAM INEG = -0.435
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
.ENDS LM358TI
*



