.SUBCKT irlb8748pbf 1 2 3
* SPICE3 MODEL WITH THERMAL RC NETWORK 
* Model generated on July 25, 11
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=2.99256 LAMBDA=0 KP=1000
+CGSO=1.95655e-05 CGDO=7.15322e-08
RS 8 3 0.00433299
D1 3 1 MD
.MODEL MD D IS=5.6658e-08 RS=0.0026978 N=1.35469 BV=30
+IBV=0.00025 EG=1.2 XTI=1.01621 TT=1e-07
+CJO=9.53372e-10 VJ=0.987007 M=0.448742 FC=0.5
RDS 3 1 1e+08
RD 9 1 0.0001
RG 2 7 8.38809
D2 4 5 MD1
.MODEL MD1 D IS=1e-32 N=50
+CJO=3.18152e-10 VJ=3.07419 M=0.3 FC=1e-08
D3 0 5 MD2
.MODEL MD2 D IS=1e-10 N=0.400002 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 9.20352e-10
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
.MODEL MD3 D IS=1e-10 N=0.400002
.ENDS irlb8748pbf


*SPICE Thermal Model Subcircuit
.SUBCKT irlb8748pbft 4 0

R_RTHERM1         4 3  1.55246
R_RTHERM2         3 2  0.00682
R_RTHERM3         2 1  0.00172
R_RTHERM4         1 0  0.43999
C_CTHERM1         4 3  0.00341
C_CTHERM2         3 2  1209.75
C_CTHERM3         2 1  4027.15
C_CTHERM4         1 0  0.00072

.ENDS irlb8748pbft

